//register file for the single cycle cpu
module register
(
input WrEn
input[31:0] Dw
);

endmodule