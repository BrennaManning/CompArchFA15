module instructionfetchunit(
	);
endmodule