module instructiondecoder(
	);
endmodule