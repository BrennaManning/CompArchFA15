module pc_register(
	input [31:0] pc_reg_in,
	output [31:0] pc_reg_out
	);

	assign pc_reg_out = pc_reg_in;

endmodule